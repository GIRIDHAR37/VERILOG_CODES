module pwm #(parameter R=8)(input clk,rst_n,
						   input [R-1:0]duty,
						   output pwm_out
						  );

	   reg [R-1:0]q_reg,q_next;

	   always @(posedge clk, negedge rst_n) begin
	   		if(~rst_n)
				q_reg<='b0;
			else
				q_reg<=q_next;
	   end

	   always @(*) begin
	   		q_next=q_reg+1;
	   end

	   assign pwm_out = (q_reg < duty);

endmodule

// output :
/*
# Time: 0, clk: 0, rst_n: 0, duty: x, pwm_out: x
# Time: 2, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 5, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 10, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 15, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 20, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 25, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 30, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 35, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 40, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 45, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 50, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 55, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 60, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 65, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 70, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 75, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 80, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 85, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 90, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 95, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 100, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 105, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 110, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 115, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 120, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 125, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 130, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 135, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 140, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 145, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 150, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 155, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 160, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 165, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 170, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 175, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 180, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 185, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 190, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 195, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 200, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 205, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 210, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 215, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 220, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 225, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 230, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 235, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 240, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 245, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 250, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 255, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 260, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 265, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 270, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 275, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 280, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 285, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 290, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 295, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 300, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 305, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 310, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 315, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 320, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 325, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 330, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 335, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 340, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 345, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 350, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 355, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 360, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 365, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 370, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 375, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 380, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 385, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 390, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 395, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 400, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 405, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 410, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 415, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 420, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 425, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 430, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 435, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 440, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 445, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 450, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 455, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 460, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 465, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 470, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 475, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 480, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 485, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 490, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 495, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 500, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 505, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 510, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 515, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 520, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 525, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 530, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 535, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 540, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 545, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 550, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 555, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 560, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 565, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 570, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 575, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 580, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 585, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 590, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 595, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 600, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 605, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 610, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 615, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 620, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 625, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 630, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 635, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 640, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 645, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 650, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 655, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 660, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 665, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 670, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 675, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 680, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 685, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 690, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 695, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 700, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 705, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 710, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 715, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 720, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 725, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 730, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 735, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 740, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 745, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 750, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 755, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 760, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 765, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 770, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 775, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 780, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 785, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 790, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 795, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 800, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 805, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 810, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 815, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 820, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 825, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 830, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 835, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 840, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 845, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 850, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 855, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 860, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 865, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 870, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 875, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 880, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 885, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 890, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 895, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 900, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 905, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 910, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 915, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 920, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 925, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 930, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 935, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 940, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 945, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 950, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 955, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 960, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 965, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 970, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 975, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 980, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 985, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 990, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 995, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1000, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1005, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1010, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1015, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1020, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1025, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1030, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1035, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1040, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1045, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1050, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1055, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1060, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1065, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1070, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1075, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1080, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1085, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1090, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1095, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1100, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1105, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1110, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1115, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1120, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1125, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1130, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1135, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1140, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1145, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1150, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1155, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1160, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1165, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1170, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1175, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1180, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1185, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1190, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1195, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1200, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1205, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1210, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1215, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1220, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1225, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1230, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1235, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1240, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1245, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1250, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1255, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1260, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1265, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1270, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1275, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1280, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1285, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1290, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1295, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1300, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1305, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1310, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1315, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1320, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1325, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1330, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1335, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1340, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1345, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1350, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1355, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1360, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1365, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1370, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1375, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1380, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1385, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1390, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1395, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1400, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1405, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1410, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1415, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1420, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1425, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1430, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1435, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1440, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1445, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1450, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1455, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1460, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1465, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1470, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1475, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1480, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1485, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1490, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1495, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1500, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1505, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1510, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1515, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1520, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1525, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1530, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1535, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1540, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1545, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1550, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1555, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1560, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1565, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1570, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1575, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1580, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1585, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1590, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1595, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1600, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1605, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1610, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1615, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1620, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1625, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1630, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1635, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1640, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1645, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1650, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1655, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1660, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1665, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1670, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1675, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1680, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1685, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1690, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1695, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1700, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1705, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1710, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1715, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1720, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1725, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1730, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1735, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1740, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1745, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1750, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1755, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1760, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1765, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1770, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1775, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1780, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1785, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1790, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1795, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1800, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1805, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1810, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1815, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1820, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1825, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1830, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1835, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1840, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1845, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1850, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1855, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1860, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1865, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1870, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1875, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1880, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1885, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1890, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1895, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1900, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1905, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1910, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1915, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1920, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1925, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1930, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1935, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1940, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1945, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1950, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1955, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1960, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1965, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1970, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1975, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1980, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1985, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1990, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 1995, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2000, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2005, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2010, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2015, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2020, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2025, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2030, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2035, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2040, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2045, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2050, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2055, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2060, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2065, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2070, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2075, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2080, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2085, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2090, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2095, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2100, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2105, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2110, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2115, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2120, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2125, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2130, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2135, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2140, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2145, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2150, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2155, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2160, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2165, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2170, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2175, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2180, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2185, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2190, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2195, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2200, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2205, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2210, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2215, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2220, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2225, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2230, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2235, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2240, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2245, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2250, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2255, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2260, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2265, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2270, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2275, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2280, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2285, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2290, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2295, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2300, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2305, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2310, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2315, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2320, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2325, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2330, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2335, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2340, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2345, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2350, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2355, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2360, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2365, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2370, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2375, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2380, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2385, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2390, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2395, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2400, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2405, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2410, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2415, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2420, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2425, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2430, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2435, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2440, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2445, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2450, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2455, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2460, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2465, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2470, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2475, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2480, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2485, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2490, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2495, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2500, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2505, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2510, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2515, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2520, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2525, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2530, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2535, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2540, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2545, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2550, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 2555, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2560, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2565, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2570, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2575, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2580, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2585, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2590, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2595, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2600, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2605, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2610, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2615, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2620, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2625, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2630, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2635, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2640, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2645, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2650, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2655, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2660, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2665, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2670, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2675, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2680, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2685, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2690, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2695, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2700, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2705, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2710, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2715, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2720, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2725, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2730, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2735, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2740, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2745, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2750, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2755, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2760, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2765, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2770, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2775, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2780, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2785, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2790, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2795, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2800, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2805, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2810, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2815, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2820, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2825, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2830, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2835, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2840, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2845, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2850, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2855, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2860, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2865, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2870, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2875, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2880, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2885, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2890, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2895, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2900, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2905, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2910, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2915, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2920, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2925, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2930, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2935, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2940, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2945, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2950, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2955, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2960, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2965, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2970, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2975, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2980, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2985, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2990, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 2995, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3000, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3005, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3010, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3015, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3020, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3025, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3030, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3035, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3040, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3045, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3050, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3055, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3060, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3065, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3070, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3075, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3080, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3085, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3090, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3095, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3100, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3105, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3110, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3115, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3120, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3125, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3130, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3135, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3140, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3145, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3150, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3155, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3160, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3165, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3170, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3175, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3180, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3185, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3190, clk: 0, rst_n: 1, duty: 64, pwm_out: 1
# Time: 3195, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3200, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3205, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3210, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3215, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3220, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3225, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3230, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3235, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3240, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3245, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3250, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3255, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3260, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3265, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3270, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3275, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3280, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3285, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3290, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3295, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3300, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3305, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3310, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3315, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3320, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3325, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3330, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3335, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3340, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3345, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3350, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3355, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3360, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3365, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3370, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3375, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3380, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3385, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3390, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3395, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3400, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3405, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3410, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3415, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3420, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3425, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3430, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3435, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3440, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3445, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3450, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3455, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3460, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3465, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3470, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3475, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3480, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3485, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3490, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3495, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3500, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3505, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3510, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3515, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3520, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3525, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3530, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3535, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3540, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3545, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3550, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3555, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3560, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3565, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3570, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3575, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3580, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3585, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3590, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3595, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3600, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3605, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3610, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3615, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3620, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3625, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3630, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3635, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3640, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3645, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3650, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3655, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3660, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3665, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3670, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3675, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3680, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3685, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3690, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3695, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3700, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3705, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3710, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3715, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3720, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3725, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3730, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3735, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3740, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3745, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3750, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3755, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3760, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3765, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3770, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3775, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3780, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3785, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3790, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3795, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3800, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3805, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3810, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3815, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3820, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3825, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3830, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3835, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3840, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3845, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3850, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3855, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3860, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3865, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3870, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3875, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3880, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3885, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3890, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3895, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3900, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3905, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3910, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3915, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3920, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3925, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3930, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3935, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3940, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3945, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3950, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3955, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3960, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3965, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3970, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3975, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3980, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3985, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3990, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 3995, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4000, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4005, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4010, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4015, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4020, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4025, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4030, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4035, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4040, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4045, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4050, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4055, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4060, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4065, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4070, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4075, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4080, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4085, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4090, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4095, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4100, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4105, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4110, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4115, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4120, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4125, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4130, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4135, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4140, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4145, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4150, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4155, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4160, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4165, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4170, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4175, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4180, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4185, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4190, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4195, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4200, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4205, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4210, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4215, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4220, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4225, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4230, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4235, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4240, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4245, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4250, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4255, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4260, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4265, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4270, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4275, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4280, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4285, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4290, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4295, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4300, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4305, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4310, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4315, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4320, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4325, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4330, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4335, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4340, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4345, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4350, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4355, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4360, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4365, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4370, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4375, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4380, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4385, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4390, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4395, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4400, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4405, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4410, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4415, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4420, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4425, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4430, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4435, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4440, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4445, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4450, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4455, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4460, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4465, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4470, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4475, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4480, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4485, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4490, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4495, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4500, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4505, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4510, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4515, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4520, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4525, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4530, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4535, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4540, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4545, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4550, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4555, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4560, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4565, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4570, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4575, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4580, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4585, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4590, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4595, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4600, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4605, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4610, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4615, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4620, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4625, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4630, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4635, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4640, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4645, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4650, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4655, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4660, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4665, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4670, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4675, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4680, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4685, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4690, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4695, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4700, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4705, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4710, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4715, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4720, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4725, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4730, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4735, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4740, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4745, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4750, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4755, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4760, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4765, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4770, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4775, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4780, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4785, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4790, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4795, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4800, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4805, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4810, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4815, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4820, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4825, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4830, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4835, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4840, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4845, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4850, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4855, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4860, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4865, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4870, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4875, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4880, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4885, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4890, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4895, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4900, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4905, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4910, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4915, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4920, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4925, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4930, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4935, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4940, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4945, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4950, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4955, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4960, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4965, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4970, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4975, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4980, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4985, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4990, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 4995, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5000, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5005, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5010, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5015, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5020, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5025, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5030, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5035, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5040, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5045, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5050, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5055, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5060, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5065, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5070, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5075, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5080, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5085, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5090, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5095, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5100, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5105, clk: 1, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5110, clk: 0, rst_n: 1, duty: 64, pwm_out: 0
# Time: 5115, clk: 1, rst_n: 1, duty: 64, pwm_out: 1
# Time: 5120, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5125, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5130, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5135, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5140, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5145, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5150, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5155, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5160, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5165, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5170, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5175, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5180, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5185, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5190, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5195, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5200, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5205, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5210, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5215, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5220, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5225, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5230, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5235, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5240, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5245, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5250, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5255, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5260, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5265, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5270, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5275, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5280, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5285, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5290, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5295, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5300, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5305, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5310, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5315, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5320, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5325, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5330, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5335, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5340, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5345, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5350, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5355, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5360, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5365, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5370, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5375, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5380, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5385, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5390, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5395, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5400, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5405, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5410, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5415, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5420, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5425, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5430, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5435, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5440, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5445, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5450, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5455, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5460, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5465, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5470, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5475, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5480, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5485, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5490, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5495, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5500, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5505, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5510, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5515, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5520, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5525, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5530, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5535, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5540, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5545, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5550, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5555, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5560, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5565, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5570, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5575, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5580, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5585, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5590, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5595, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5600, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5605, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5610, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5615, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5620, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5625, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5630, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5635, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5640, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5645, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5650, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5655, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5660, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5665, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5670, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5675, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5680, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5685, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5690, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5695, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5700, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5705, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5710, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5715, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5720, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5725, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5730, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5735, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5740, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5745, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5750, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5755, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5760, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5765, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5770, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5775, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5780, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5785, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5790, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5795, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5800, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5805, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5810, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5815, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5820, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5825, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5830, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5835, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5840, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5845, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5850, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5855, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5860, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5865, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5870, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5875, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5880, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5885, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5890, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5895, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5900, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5905, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5910, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5915, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5920, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5925, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5930, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5935, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5940, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5945, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5950, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5955, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5960, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5965, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5970, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5975, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5980, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5985, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5990, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 5995, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6000, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6005, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6010, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6015, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6020, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6025, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6030, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6035, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6040, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6045, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6050, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6055, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6060, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6065, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6070, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6075, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6080, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6085, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6090, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6095, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6100, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6105, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6110, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6115, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6120, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6125, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6130, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6135, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6140, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6145, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6150, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6155, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6160, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6165, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6170, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6175, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6180, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6185, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6190, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6195, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6200, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6205, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6210, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6215, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6220, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6225, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6230, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6235, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6240, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6245, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6250, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6255, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6260, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6265, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6270, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6275, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6280, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6285, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6290, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6295, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6300, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6305, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6310, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6315, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6320, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6325, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6330, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6335, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6340, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6345, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6350, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6355, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6360, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6365, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6370, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6375, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6380, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6385, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6390, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 6395, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6400, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6405, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6410, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6415, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6420, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6425, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6430, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6435, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6440, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6445, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6450, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6455, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6460, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6465, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6470, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6475, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6480, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6485, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6490, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6495, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6500, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6505, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6510, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6515, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6520, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6525, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6530, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6535, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6540, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6545, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6550, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6555, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6560, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6565, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6570, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6575, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6580, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6585, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6590, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6595, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6600, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6605, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6610, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6615, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6620, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6625, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6630, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6635, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6640, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6645, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6650, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6655, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6660, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6665, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6670, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6675, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6680, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6685, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6690, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6695, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6700, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6705, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6710, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6715, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6720, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6725, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6730, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6735, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6740, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6745, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6750, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6755, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6760, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6765, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6770, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6775, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6780, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6785, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6790, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6795, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6800, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6805, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6810, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6815, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6820, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6825, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6830, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6835, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6840, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6845, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6850, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6855, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6860, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6865, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6870, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6875, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6880, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6885, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6890, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6895, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6900, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6905, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6910, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6915, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6920, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6925, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6930, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6935, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6940, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6945, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6950, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6955, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6960, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6965, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6970, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6975, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6980, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6985, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6990, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 6995, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7000, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7005, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7010, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7015, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7020, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7025, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7030, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7035, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7040, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7045, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7050, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7055, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7060, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7065, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7070, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7075, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7080, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7085, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7090, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7095, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7100, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7105, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7110, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7115, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7120, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7125, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7130, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7135, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7140, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7145, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7150, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7155, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7160, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7165, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7170, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7175, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7180, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7185, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7190, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7195, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7200, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7205, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7210, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7215, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7220, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7225, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7230, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7235, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7240, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7245, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7250, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7255, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7260, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7265, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7270, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7275, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7280, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7285, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7290, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7295, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7300, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7305, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7310, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7315, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7320, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7325, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7330, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7335, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7340, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7345, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7350, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7355, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7360, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7365, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7370, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7375, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7380, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7385, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7390, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7395, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7400, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7405, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7410, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7415, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7420, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7425, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7430, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7435, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7440, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7445, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7450, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7455, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7460, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7465, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7470, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7475, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7480, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7485, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7490, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7495, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7500, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7505, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7510, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7515, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7520, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7525, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7530, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7535, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7540, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7545, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7550, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7555, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7560, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7565, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7570, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7575, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7580, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7585, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7590, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7595, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7600, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7605, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7610, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7615, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7620, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7625, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7630, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7635, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7640, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7645, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7650, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7655, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7660, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7665, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7670, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 7675, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7680, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7685, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7690, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7695, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7700, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7705, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7710, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7715, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7720, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7725, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7730, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7735, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7740, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7745, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7750, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7755, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7760, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7765, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7770, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7775, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7780, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7785, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7790, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7795, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7800, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7805, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7810, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7815, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7820, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7825, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7830, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7835, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7840, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7845, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7850, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7855, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7860, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7865, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7870, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7875, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7880, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7885, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7890, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7895, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7900, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7905, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7910, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7915, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7920, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7925, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7930, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7935, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7940, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7945, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7950, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7955, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7960, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7965, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7970, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7975, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7980, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7985, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7990, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 7995, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8000, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8005, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8010, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8015, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8020, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8025, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8030, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8035, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8040, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8045, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8050, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8055, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8060, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8065, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8070, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8075, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8080, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8085, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8090, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8095, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8100, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8105, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8110, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8115, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8120, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8125, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8130, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8135, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8140, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8145, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8150, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8155, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8160, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8165, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8170, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8175, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8180, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8185, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8190, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8195, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8200, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8205, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8210, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8215, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8220, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8225, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8230, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8235, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8240, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8245, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8250, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8255, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8260, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8265, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8270, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8275, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8280, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8285, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8290, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8295, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8300, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8305, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8310, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8315, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8320, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8325, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8330, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8335, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8340, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8345, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8350, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8355, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8360, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8365, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8370, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8375, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8380, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8385, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8390, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8395, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8400, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8405, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8410, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8415, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8420, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8425, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8430, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8435, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8440, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8445, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8450, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8455, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8460, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8465, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8470, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8475, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8480, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8485, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8490, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8495, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8500, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8505, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8510, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8515, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8520, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8525, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8530, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8535, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8540, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8545, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8550, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8555, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8560, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8565, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8570, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8575, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8580, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8585, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8590, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8595, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8600, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8605, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8610, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8615, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8620, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8625, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8630, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8635, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8640, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8645, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8650, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8655, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8660, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8665, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8670, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8675, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8680, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8685, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8690, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8695, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8700, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8705, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8710, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8715, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8720, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8725, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8730, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8735, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8740, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8745, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8750, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8755, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8760, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8765, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8770, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8775, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8780, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8785, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8790, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8795, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8800, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8805, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8810, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8815, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8820, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8825, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8830, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8835, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8840, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8845, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8850, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8855, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8860, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8865, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8870, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8875, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8880, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8885, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8890, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8895, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8900, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8905, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8910, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8915, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8920, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8925, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8930, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8935, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8940, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8945, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8950, clk: 0, rst_n: 1, duty: 128, pwm_out: 1
# Time: 8955, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8960, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8965, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8970, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8975, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8980, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8985, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8990, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 8995, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9000, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9005, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9010, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9015, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9020, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9025, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9030, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9035, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9040, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9045, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9050, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9055, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9060, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9065, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9070, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9075, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9080, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9085, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9090, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9095, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9100, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9105, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9110, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9115, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9120, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9125, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9130, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9135, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9140, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9145, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9150, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9155, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9160, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9165, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9170, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9175, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9180, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9185, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9190, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9195, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9200, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9205, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9210, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9215, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9220, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9225, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9230, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9235, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9240, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9245, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9250, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9255, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9260, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9265, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9270, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9275, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9280, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9285, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9290, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9295, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9300, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9305, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9310, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9315, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9320, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9325, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9330, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9335, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9340, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9345, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9350, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9355, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9360, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9365, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9370, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9375, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9380, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9385, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9390, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9395, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9400, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9405, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9410, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9415, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9420, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9425, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9430, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9435, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9440, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9445, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9450, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9455, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9460, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9465, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9470, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9475, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9480, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9485, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9490, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9495, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9500, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9505, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9510, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9515, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9520, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9525, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9530, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9535, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9540, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9545, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9550, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9555, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9560, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9565, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9570, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9575, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9580, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9585, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9590, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9595, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9600, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9605, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9610, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9615, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9620, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9625, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9630, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9635, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9640, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9645, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9650, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9655, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9660, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9665, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9670, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9675, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9680, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9685, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9690, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9695, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9700, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9705, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9710, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9715, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9720, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9725, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9730, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9735, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9740, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9745, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9750, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9755, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9760, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9765, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9770, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9775, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9780, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9785, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9790, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9795, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9800, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9805, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9810, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9815, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9820, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9825, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9830, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9835, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9840, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9845, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9850, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9855, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9860, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9865, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9870, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9875, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9880, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9885, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9890, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9895, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9900, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9905, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9910, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9915, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9920, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9925, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9930, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9935, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9940, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9945, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9950, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9955, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9960, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9965, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9970, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9975, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9980, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9985, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9990, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 9995, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10000, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10005, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10010, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10015, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10020, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10025, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10030, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10035, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10040, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10045, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10050, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10055, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10060, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10065, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10070, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10075, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10080, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10085, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10090, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10095, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10100, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10105, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10110, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10115, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10120, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10125, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10130, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10135, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10140, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10145, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10150, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10155, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10160, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10165, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10170, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10175, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10180, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10185, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10190, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10195, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10200, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10205, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10210, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10215, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10220, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10225, clk: 1, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10230, clk: 0, rst_n: 1, duty: 128, pwm_out: 0
# Time: 10235, clk: 1, rst_n: 1, duty: 128, pwm_out: 1
# Time: 10240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10275, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10280, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10285, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10290, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10295, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10300, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10305, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10310, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10315, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10320, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10325, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10330, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10335, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10340, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10345, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10350, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10715, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10720, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10725, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10730, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10735, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10740, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10745, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10750, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10755, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10760, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10765, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10770, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10775, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10780, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10785, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10790, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 10995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11155, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11160, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11165, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11170, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11175, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11180, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11185, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11190, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11195, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11200, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11205, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11210, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11215, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11220, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11225, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11230, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11235, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11275, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11280, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11285, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11290, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11295, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11300, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11305, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11310, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11315, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11320, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11325, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11330, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11335, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11340, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11345, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11350, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11715, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11720, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11725, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11730, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11735, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11740, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11745, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11750, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11755, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11760, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11765, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11770, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11775, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11780, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11785, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11790, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 11995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12155, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12160, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12165, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12170, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12175, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12180, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12185, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12190, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12195, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12200, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12205, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12210, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12215, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12220, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12225, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12230, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12235, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12240, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12245, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12250, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12255, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12260, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12265, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12270, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12275, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12280, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12285, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12290, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12295, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12300, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12305, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12310, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12315, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12320, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12325, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12330, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12335, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12340, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12345, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12350, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12355, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12360, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12365, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12370, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12375, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12380, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12385, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12390, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12395, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12400, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12405, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12410, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12415, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12420, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12425, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12430, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12435, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12440, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12445, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12450, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12455, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12460, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12465, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12470, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12475, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12480, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12485, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12490, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12495, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12500, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12505, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12510, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12515, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12520, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12525, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12530, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12535, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12540, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12545, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12550, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12555, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12560, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12565, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12570, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12575, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12580, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12585, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12590, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12595, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12600, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12605, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12610, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12615, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12620, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12625, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12630, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12635, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12640, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12645, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12650, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12655, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12660, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12665, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12670, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12675, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12680, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12685, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12690, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12695, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12700, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12705, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12710, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12715, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12720, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12725, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12730, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12735, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12740, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12745, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12750, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12755, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12760, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12765, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12770, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12775, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12780, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12785, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12790, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 12795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 12995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13155, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13160, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13165, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13170, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13175, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13180, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13185, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13190, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13195, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13200, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13205, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13210, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13215, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13220, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13225, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13230, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13235, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13275, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13280, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13285, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13290, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13295, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13300, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13305, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13310, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13315, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13320, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13325, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13330, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13335, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13340, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13345, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13350, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13715, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13720, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13725, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13730, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13735, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13740, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13745, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13750, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13755, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13760, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13765, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13770, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13775, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13780, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13785, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13790, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 13995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14155, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14160, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14165, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14170, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14175, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14180, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14185, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14190, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14195, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14200, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14205, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14210, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14215, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14220, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14225, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14230, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14235, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14275, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14280, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14285, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14290, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14295, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14300, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14305, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14310, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14315, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14320, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14325, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14330, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14335, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14340, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14345, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14350, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 14715, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14720, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14725, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14730, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14735, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14740, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14745, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14750, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14755, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14760, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14765, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14770, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14775, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14780, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14785, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14790, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14795, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14800, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14805, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14810, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14815, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14820, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14825, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14830, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14835, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14840, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14845, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14850, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14855, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14860, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14865, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14870, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14875, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14880, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14885, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14890, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14895, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14900, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14905, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14910, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14915, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14920, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14925, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14930, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14935, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14940, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14945, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14950, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14955, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14960, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14965, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14970, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14975, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14980, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14985, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14990, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 14995, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15000, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15005, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15010, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15015, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15020, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15025, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15030, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15035, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15040, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15045, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15050, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15055, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15060, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15065, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15070, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15075, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15080, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15085, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15090, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15095, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15100, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15105, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15110, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15115, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15120, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15125, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15130, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15135, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15140, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15145, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15150, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15155, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15160, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15165, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15170, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15175, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15180, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15185, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15190, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15195, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15200, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15205, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15210, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15215, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15220, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15225, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15230, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15235, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15240, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15245, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15250, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15255, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15260, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15265, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15270, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15275, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15280, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15285, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15290, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15295, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15300, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15305, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15310, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15315, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15320, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15325, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15330, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15335, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15340, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15345, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15350, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 15355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15715, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15720, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15725, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15730, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15735, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15740, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15745, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15750, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15755, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15760, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15765, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15770, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15775, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15780, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15785, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15790, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 15995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16155, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16160, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16165, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16170, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16175, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16180, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16185, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16190, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16195, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16200, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16205, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16210, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16215, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16220, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16225, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16230, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16235, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16275, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16280, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16285, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16290, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16295, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16300, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16305, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16310, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16315, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16320, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16325, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16330, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16335, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16340, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16345, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16350, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16355, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16360, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16365, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16370, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16375, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16380, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16385, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16390, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16395, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16400, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16405, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16410, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16415, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16420, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16425, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16430, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16435, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16440, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16445, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16450, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16455, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16460, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16465, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16470, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16475, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16480, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16485, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16490, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16495, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16500, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16505, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16510, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16515, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16520, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16525, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16530, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16535, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16540, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16545, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16550, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16555, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16560, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16565, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16570, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16575, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16580, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16585, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16590, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16595, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16600, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16605, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16610, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16615, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16620, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16625, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16630, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16635, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16640, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16645, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16650, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16655, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16660, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16665, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16670, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16675, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16680, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16685, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16690, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16695, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16700, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16705, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16710, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16715, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16720, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16725, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16730, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16735, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16740, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16745, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16750, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16755, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16760, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16765, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16770, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16775, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16780, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16785, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16790, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16795, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16800, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16805, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16810, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16815, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16820, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16825, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16830, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16835, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16840, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16845, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16850, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16855, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16860, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16865, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16870, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16875, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16880, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16885, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16890, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16895, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16900, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16905, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16910, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16920, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16925, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16930, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16935, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16940, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16945, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16950, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16955, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16960, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16965, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16970, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16975, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16980, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16985, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16990, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 16995, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17000, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17005, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17010, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17015, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17020, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17025, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17030, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17035, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17040, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17045, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17050, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17055, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17060, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17065, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17070, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17075, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17080, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17085, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17090, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17095, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17100, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17105, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17110, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17115, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17120, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17125, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17130, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17135, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17140, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17145, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17150, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17155, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17160, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17165, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17170, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17175, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17180, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17185, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17190, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17195, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17200, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17205, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17210, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17215, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17220, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17225, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17230, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17235, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17240, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17245, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17250, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17255, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17260, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17265, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17270, clk: 0, rst_n: 1, duty: 192, pwm_out: 1
# Time: 17275, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17280, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17285, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17290, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17295, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17300, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17305, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17310, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17315, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17320, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17325, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17330, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17335, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17340, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17345, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17350, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17355, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17360, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17365, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17370, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17375, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17380, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17385, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17390, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17395, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17400, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17405, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17410, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17415, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17420, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17425, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17430, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17435, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17440, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17445, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17450, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17455, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17460, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17465, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17470, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17475, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17480, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17485, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17490, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17495, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17500, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17505, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17510, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17515, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17520, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17525, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17530, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17535, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17540, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17545, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17550, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17555, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17560, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17565, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17570, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17575, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17580, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17585, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17590, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17595, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17600, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17605, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17610, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17615, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17620, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17625, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17630, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17635, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17640, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17645, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17650, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17655, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17660, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17665, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17670, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17675, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17680, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17685, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17690, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17695, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17700, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17705, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17710, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17715, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17720, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17725, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17730, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17735, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17740, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17745, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17750, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17755, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17760, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17765, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17770, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17775, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17780, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17785, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17790, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17795, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17800, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17805, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17810, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17815, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17820, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17825, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17830, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17835, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17840, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17845, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17850, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17855, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17860, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17865, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17870, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17875, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17880, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17885, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17890, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17895, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17900, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17905, clk: 1, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17910, clk: 0, rst_n: 1, duty: 192, pwm_out: 0
# Time: 17915, clk: 1, rst_n: 1, duty: 192, pwm_out: 1
# ** Note: $stop    : pwm_tb.v(18)
#    Time: 17920 ps  Iteration: 0  Instance: /pwm_tb
*/
